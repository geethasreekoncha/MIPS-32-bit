module pipe_MIPS32 (clk1, clk2);
input clk1, clk2;
reg [31:0] PC, IF_ID_IR, IF_ID_NPC;
reg [31:0] ID_EX_IR, ID_EX_NPC, ID_EX_B, ID_EX_Imm;
reg [2:0] ID_EX_type, EX_MEM_type, MEM_WB_type;
reg EX_MEM_cond;
reg [31:0] MEM_WB_IR, MEM_WB_ALUOut, MEM_WB_LMD;
reg [31:0] Reg [0:31];
reg [31:0] Mem [0:1023];
parameter ADD=6'b000000, SUB=6'b000001, AND=6'b000010, OR=6'b000011, SLT=6'b000100, MUL=6'b000101, HLT=6'b111111, LW=6'b001000, SW=6'b001001, ADDI=6'b001010, SUBI=6'b001011, SLTI=6'b001100,
BNEQZ=6'b001101, BEQZ=6'b001110;
parameter RR_ALU=3'b000, RM_ALU=3'b001, LOAD=3'b010, STORE=3'b011, BRANCH=3'b100, HALT=3'b101;
reg HALTED;
reg TAKEN_BRANCH;
//IF stage
always @(posedge clk1)
if(HALTED==0)
begin
if (((EX_MEM_IR[31:26] == BEQZ) && (EX_MEM_cond ==1)) || ((EX_MEM_IR[31:26]== BNEQZ) && (EX_MEM_cond ==0)))
beginIF_ID_IR <= #2 Mem[EX_MEM_ALUOut];
TAKEN_BRANCH <= #2 1'b1;
IF_ID_NPC <= #2 EX_MEM_ALUOut +1;
PC <= #2 EX_MEM_ALUOut +1;
end
else
begin
IF_ID_IR <= #2 Mem[PC];
IF_ID_NPC <= PC +1;
PC <= #2 PC +1;
end
end

//ID stage
always @(posedge clk2)
if(HALTED == 0)
begin
if(IF_ID_IR[25:21] == 5'b00000) ID_EX_A <=0;
else ID_EX_A <= #2 Reg[IF_ID_IR[25:21]];

if(IF_ID_IR[20:16] == 5'b00000) ID_EX_B <=0;
else ID_EX_B <= #2 Reg[IF_IR[20:16]];

ID_EX_NPC <= #2 IF_ID_NPC;
ID_EX_IR <= #2 IF_ID_IR;
ID_EX_Imm <= #2 {{16{IF_ID_IR[15]}}, {IF_ID_IR[15:0]}};
